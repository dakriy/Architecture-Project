alu.
